module main

fn main(){
	println("Not available...")
}