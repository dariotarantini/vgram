module hygram

import http
import json


// main struct
struct Telegram {
    Token string
}
