module vgram
// getUpdates
pub struct NewGetUpdates {
pub:
    offset int
    limit int
    timeout int
    allowed_updates []string
}
// sendMessage
pub struct NewSendMessage {
pub:
    chat_id string
    text string
    parse_mode string
    disable_web_page_preview bool
    disable_notification bool
    reply_to_message_id int
    reply_markup string
}
// forwardMessage
pub struct NewForwardMessage {
pub:
    chat_id string
	from_chat_id string
	disable_notification bool
	message_id int
}
// sendPhoto
pub struct NewSendPhoto {
pub:
    chat_id string
	photo string
    caption string
    parse_mode string
    disable_web_page_preview bool
    disable_notification bool
    reply_to_message_id int
    reply_markup string
}
// sendAudio
pub struct NewSendAudio {
pub:
    chat_id string
	audio string
    caption string
    parse_mode string
	performer string
	title string
	thumb string
    disable_notification bool
    reply_to_message_id int
    reply_markup string
}
// sendDocument
pub struct NewSendDocument {
pub:
    chat_id string
	document string
    caption string
    parse_mode string
	thumb string
    disable_notification bool
    reply_to_message_id int
    reply_markup string
}
// sendVideo
pub struct NewSendVideo {
pub:
    chat_id string
	video string
	duration int
	width int
	height int
	supports_streaming bool
    caption string
    parse_mode string
	thumb string
    disable_notification bool
    reply_to_message_id int
    reply_markup string
}
// sendAnimation
pub struct NewSendAnimation {
pub:
    chat_id string
	animation string
	duration int
	width int
	height int
    caption string
    parse_mode string
	thumb string
    disable_notification bool
    reply_to_message_id int
    reply_markup string
}
// sendVoice
pub struct NewSendVoice {
pub:
    chat_id string
	voice string
	duration int
    caption string
    parse_mode string
	thumb string
    disable_notification bool
    reply_to_message_id int
    reply_markup string
}
// sendVideoNote
pub struct NewSendVideoNote {
pub:
    chat_id string
	video_note string
	duration int
	length int
    caption string
    parse_mode string
	thumb string
    disable_notification bool
    reply_to_message_id int
    reply_markup string
}
// sendMediaGroup
pub struct NewSendMediaGroup {
pub:
    chat_id string
	media string // json of []InputMedia (not implemented)
    disable_notification bool
    reply_to_message_id int
    reply_markup string
}
// sendLocation
pub struct NewSendLocation {
pub:
    chat_id string
	latitude f32
	longitude f32
	live_period int
    disable_notification bool
    reply_to_message_id int
    reply_markup string
}
// editMessageLiveLocation
pub struct NewEditMessageLiveLocation {
pub:
    chat_id string
	message_id int
	inline_message_id string
	latitude f32
    longitude f32
    reply_markup string
}
// stopMessageLiveLocation
pub struct NewStopMessageLiveLocation {
pub:
    chat_id string
	message_id int
	inline_message_id string
    reply_markup string
}
// sendVenue
pub struct NewSendVenue {
pub:
    chat_id string
	latitude f32
    longitude  f32
    title string
    address string
    foursquare_id string
    foursquare_type string
    disable_notification bool
    reply_to_message_id int
    reply_markup string
}
// sendContact
pub struct NewSendContact {
pub:
    chat_id string
    phone_number string
    first_name string
    last_name string
    vcard string
    disable_notification bool
    reply_to_message_id int
    reply_markup string
}
// sendPoll
pub struct NewSendPoll {
pub:
    chat_id string
    question string
    options []string
    disable_notification bool
    reply_to_message_id int
    reply_markup string
}
// sendChatAction
pub struct NewSendChatAction {
pub:
    chat_id string
    action string
}
// getUserProfilePhotos
pub struct NewGetUserProfilePhotos {
pub:
    user_id int
    offset int
    limit int
}
// getFile
pub struct NewGetFile {
pub:
    file_id string
}
pub struct NewAnswerInlineQuery {
pub:
    inline_query_id string
    results string  // json of []InlineQueryResult (not implemented)
    cache_time int
    is_personal int
    next_offset string
    switch_pm_text string
    switch_pm_parameter string
}